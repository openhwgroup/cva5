/*
 * Copyright © 2019-2023 Yuhui Gao, Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Yuhui Gao <yuhuig@sfu.ca>
 */

module parallel_OR
#(
    parameter WIDTH
)(
    input logic [I_WIDTH-1:0] i_data,
    output logic [WIDTH-1:0] o_data
);
    localparam I_WIDTH = WIDTH*6;

    genvar i;
    generate
        for (i = 0; i < WIDTH; i++) begin
            assign o_data[i] = |i_data[6*i+:6];
        end
    endgenerate

endmodule
