/*
 * Copyright © 2020 Eric Matthews,  Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Yuhui Gao <yuhuig@sfu.ca>
 */

module fp_register_file

    import taiga_config::*;
    import riscv_types::*;
    import taiga_types::*;
     # (
        parameter cpu_config_t CONFIG = EXAMPLE_CONFIG
    )
    (
        input logic clk,
        input logic rst,
        input gc_outputs_t gc,

        //decode write interface
        input phys_addr_t decode_phys_rs_addr [FP_REGFILE_READ_PORTS],
        //input logic [$clog2(CONFIG.FP.FP_NUM_WB_GROUPS)-1:0] decode_rs_wb_group [FP_REGFILE_READ_PORTS],
        input logic decode_rs_wb_group [FP_REGFILE_READ_PORTS],
        input phys_addr_t decode_phys_rd_addr,
        input logic decode_advance,
        input logic decode_uses_rd,

        //Issue interface
        fp_register_file_issue_interface.register_file rf_issue,

        //Writeback
        input fp_commit_packet_t commit [FP_NUM_WB_GROUPS]
    );
    typedef logic [FLEN-1:0] rs_data_set_t [FP_REGFILE_READ_PORTS];
    rs_data_set_t rs_data_set [FP_NUM_WB_GROUPS];

    logic decode_inuse [FP_REGFILE_READ_PORTS];
    logic decode_inuse_r [FP_REGFILE_READ_PORTS];

    genvar i;
    ////////////////////////////////////////////////////
    //Implementation

    ////////////////////////////////////////////////////
    //Phys register inuse
    //toggle ports: decode advance, single-cycle/fetch_flush, multi-cycle commit
    //read ports: rs-decode, rs-issue

    toggle_memory_set # (
        .DEPTH (64),
        .NUM_WRITE_PORTS (3),
        .NUM_READ_PORTS (FP_REGFILE_READ_PORTS*2),
        .WRITE_INDEX_FOR_RESET (0),
        .READ_INDEX_FOR_RESET (0)
    ) id_inuse_toggle_mem_set
    (
        .clk (clk),
        .rst (rst),
        .init_clear (gc.init_clear),
        .toggle ('{
            (decode_advance & decode_uses_rd & ~gc.fetch_flush),
            rf_issue.single_cycle_or_flush,
            commit[0].valid
        }),
        .toggle_addr ('{
            decode_phys_rd_addr, 
            rf_issue.phys_rd_addr, 
            commit[0].phys_addr
        }),
        .read_addr ('{
            decode_phys_rs_addr[RS1], 
            decode_phys_rs_addr[RS2], 
            decode_phys_rs_addr[RS3], 
            rf_issue.phys_rs_addr[RS1], 
            rf_issue.phys_rs_addr[RS2],
            rf_issue.phys_rs_addr[RS3]
        }),
        .in_use ('{
            decode_inuse[RS1],
            decode_inuse[RS2],
            decode_inuse[RS3],
            rf_issue.inuse[RS1],
            rf_issue.inuse[RS2],
            rf_issue.inuse[RS3]
        })
    );
    always_ff @ (posedge clk) begin
        if (decode_advance)
            decode_inuse_r <= decode_inuse;
    end
    ////////////////////////////////////////////////////
    //Register Banks
    //Implemented in seperate module as there is not universal tool support for inferring
    //arrays of memory blocks.
    generate for (i = 0; i < FP_NUM_WB_GROUPS; i++) begin : register_file_gen
        fp_register_bank #(.NUM_READ_PORTS(FP_REGFILE_READ_PORTS))
        reg_group (
            .clk, .rst,
            .write_addr(commit[i].phys_addr),
            .new_data(commit[i].data),
            .commit(commit[i].valid),
            .read_addr(decode_phys_rs_addr),
            .data(rs_data_set[i])
        );
    end endgenerate

    ////////////////////////////////////////////////////
    //Register File Muxing
    //logic [$clog2(CONFIG.FP.FP_NUM_WB_GROUPS)-1:0] rs_wb_group [FP_REGFILE_READ_PORTS];
    logic rs_wb_group [FP_REGFILE_READ_PORTS];
    logic bypass [FP_REGFILE_READ_PORTS];
    assign rs_wb_group = decode_advance ? decode_rs_wb_group : rf_issue.rs_wb_group;
    assign bypass = decode_advance ? decode_inuse : decode_inuse_r;

    always_ff @ (posedge clk) begin
       for (int i = 0; i < FP_REGFILE_READ_PORTS; i++) begin
           if (decode_advance | rf_issue.inuse[i])
               rf_issue.data[i] <= bypass[i] ? commit[rs_wb_group[i]].data : rs_data_set[rs_wb_group[i]][i];
       end
   end

    ////////////////////////////////////////////////////
    //End of Implementation
    ////////////////////////////////////////////////////

    ////////////////////////////////////////////////////
    //Assertions
    //for (genvar i = 0; i < FP_NUM_WB_GROUPS; i++) begin : write_to_rd_zero_assertion
        //assert property (@(posedge clk) disable iff (rst) (commit[i].valid) |-> (commit[i].phys_addr != 0)) else $error("write to register zero");
    //end

endmodule
