/*
 * Copyright © 2019-2023 Yuhui Gao, Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Yuhui Gao <yuhuig@sfu.ca>
 */

//Misc. floating-point units that write-back to integer register file
//Sharing 1 write-back port
//FCMP, FCLASS, F2I
module fp_wb2int_misc
    import taiga_config::*;
    import riscv_types::*;
    import taiga_types::*;
    import fpu_types::*;

(
    input logic clk,
    unit_issue_interface.unit issue,
    input fp_wb2int_misc_inputs_t fp_wb2int_misc_inputs,
    unit_writeback_interface.unit wb
);

    fp_mv_f2i_inputs_t fp_mv_f2i_inputs;
    fp_f2i_inputs_t fp_f2i_inputs;
    fp_cmp_inputs_t fp_cmp_inputs;
    fp_class_inputs_t fp_class_inputs;
    unit_issue_interface mv_f2i_issue();
    unit_issue_interface f2i_issue();
    unit_issue_interface cmp_issue();
    unit_issue_interface class_issue();
    unit_writeback_interface mv_f2i_wb();
    unit_writeback_interface f2i_wb();
    unit_writeback_interface cmp_wb();
    unit_writeback_interface class_wb();
    logic [3:0] instruction;
    logic advance;

    ////////////////////////////////////////////////////
    //construct inputs for each unit
    assign fp_mv_f2i_inputs = fp_wb2int_misc_inputs.fp_mv_f2i_inputs;

    assign fp_f2i_inputs = fp_wb2int_misc_inputs.fp_f2i_inputs;

    assign fp_cmp_inputs = fp_wb2int_misc_inputs.fp_cmp_inputs;

    assign fp_class_inputs = fp_wb2int_misc_inputs.fp_class_inputs;

    ////////////////////////////////////////////////////
    //Issue Interfaces
    always_comb begin
        //Don't need to AND new_request with the current instruction, as the output mux handles result selection. Keeping for now for sanity check
        mv_f2i_issue.new_request = issue.new_request & fp_wb2int_misc_inputs.instruction[3];
        mv_f2i_issue.id = issue.id;
        
        f2i_issue.new_request = issue.new_request & fp_wb2int_misc_inputs.instruction[2];
        f2i_issue.id = issue.id;

        cmp_issue.new_request = issue.new_request & fp_wb2int_misc_inputs.instruction[1];
        cmp_issue.id = issue.id;

        class_issue.new_request = issue.new_request & fp_wb2int_misc_inputs.instruction[0];
        class_issue.id = issue.id;
    end

    ////////////////////////////////////////////////////
    //Mv F2I
    fp_mv_f2i fp_mv_f2i_inst(
        .clk (clk),
        .advance (advance),
        .issue (mv_f2i_issue),
        .fp_mv_f2i_inputs (fp_mv_f2i_inputs),
        .wb (mv_f2i_wb)
    );

    ////////////////////////////////////////////////////
    //F2I
    fp_f2i fp_f2i_inst(
        .clk (clk),
        .advance (advance),
        .issue (f2i_issue),
        .fp_f2i_inputs (fp_f2i_inputs),
        .wb (f2i_wb)
    );

    ////////////////////////////////////////////////////
    //FCMP
    fp_cmp fp_cmp_inst(
        .clk (clk),
        .advance (advance),
        .issue (cmp_issue),
        .fp_cmp_inputs (fp_cmp_inputs),
        .wb (cmp_wb)
    );

    ////////////////////////////////////////////////////
    //FCLASS
    fp_class fp_class_inst(
        .clk (clk),
        .advance (advance),
        .issue (class_issue),
        .fp_class_inputs (fp_class_inputs),
        .wb (class_wb)
    );

    ////////////////////////////////////////////////////
    //Control Signal
    //TODO: separate the two stages'd advance signal
    assign advance = wb.ack | ~wb.done;
    assign issue.ready = advance;

    ////////////////////////////////////////////////////
    //Registers
    always_ff @ (posedge clk) begin
        if (advance) begin
            instruction <= fp_wb2int_misc_inputs.instruction;
        end
    end

    ////////////////////////////////////////////////////
    //Output
    always_comb begin
        case(instruction)
            4'b1000: begin
                wb.done = mv_f2i_wb.done;
                wb.id = mv_f2i_wb.id;
                wb.rd = mv_f2i_wb.rd;
                wb.fflags = mv_f2i_wb.fflags;
            end
            4'b0100: begin
                wb.done = f2i_wb.done;
                wb.id = f2i_wb.id;
                wb.rd = f2i_wb.rd;
                wb.fflags = f2i_wb.fflags;
            end
            4'b0010: begin
                wb.done = cmp_wb.done;
                wb.id = cmp_wb.id;
                wb.rd = cmp_wb.rd;
                wb.fflags = cmp_wb.fflags;
            end
            default: begin
                wb.done = class_wb.done;
                wb.id = class_wb.id;
                wb.rd = class_wb.rd;
                wb.fflags = class_wb.fflags;
            end
        endcase
    end
endmodule
