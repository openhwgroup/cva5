/*
 * Copyright © 2019-2023 Yuhui Gao, Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Yuhui Gao <yuhuig@sfu.ca>
 */

module  fp_illegal_instruction_checker
    import taiga_config::*;
    import riscv_types::*;
(
    input logic [31:0] instruction,
    output logic need_int_data,
    output logic write_int_data,
    output logic need_float_data,
    output logic write_float_data,
    output logic float_instruction,
    output logic accumulating_csrs
);

    ////////////////////////////////////////////////////
    //FP instructions
    //Single Precision
    localparam [31:0] FLW       = 32'b?????????????????010?????0000111;
    localparam [31:0] FSW       = 32'b?????????????????010?????0100111;
    localparam [31:0] FMADD_S   = 32'b?????00??????????????????1000011;
    localparam [31:0] FMSUB_S   = 32'b?????00??????????????????1000111;
    localparam [31:0] FNMSUB_S  = 32'b?????00??????????????????1001011;
    localparam [31:0] FNMADD_S  = 32'b?????00??????????????????1001111;
    localparam [31:0] FADD_S    = 32'b0000000??????????????????1010011;
    localparam [31:0] FSUB_S    = 32'b0000100??????????????????1010011;
    localparam [31:0] FMUL_S    = 32'b0001000??????????????????1010011;
    localparam [31:0] FDIV_S    = 32'b0001100??????????????????1010011;
    localparam [31:0] FSQRT_S   = 32'b010110000000?????????????1010011;
    localparam [31:0] FSGNJ_S   = 32'b0010000??????????000?????1010011;
    localparam [31:0] FSGNJN_S  = 32'b0010000??????????001?????1010011;
    localparam [31:0] FSGNJX_S  = 32'b0010000??????????010?????1010011;
    localparam [31:0] FMIN_S    = 32'b0010100??????????000?????1010011;
    localparam [31:0] FMAX_S    = 32'b0010100??????????001?????1010011;
    localparam [31:0] FCVT_W_S  = 32'b110000000000?????????????1010011;
    localparam [31:0] FCVT_WU_S = 32'b110000000001?????????????1010011;
    localparam [31:0] FCVT_S_W  = 32'b110100000000?????????????1010011;
    localparam [31:0] FCVT_S_WU = 32'b110100000001?????????????1010011;
    localparam [31:0] FMV_X_W   = 32'b111000000000?????000?????1010011;
    localparam [31:0] FMV_W_X   = 32'b111100000000?????000?????1010011;
    localparam [31:0] FEQ_S     = 32'b1010000??????????010?????1010011;
    localparam [31:0] FLT_S     = 32'b1010000??????????001?????1010011;
    localparam [31:0] FLE_S     = 32'b1010000??????????000?????1010011;
    localparam [31:0] FLASS_S   = 32'b111000000000?????001?????1010011;
    //Double Precision
    localparam [31:0] FLD       = 32'b?????????????????011?????0000111;
    localparam [31:0] FSD       = 32'b?????????????????011?????0100111;
    localparam [31:0] FMADD_D   = 32'b?????01??????????????????1000011;
    localparam [31:0] FMSUB_D   = 32'b?????01??????????????????1000111;
    localparam [31:0] FNMSUB_D  = 32'b?????01??????????????????1001011;
    localparam [31:0] FNMADD_D  = 32'b?????01??????????????????1001111;
    localparam [31:0] FADD_D    = 32'b0000001??????????????????1010011;
    localparam [31:0] FSUB_D    = 32'b0000101??????????????????1010011;
    localparam [31:0] FMUL_D    = 32'b0001001??????????????????1010011;
    localparam [31:0] FDIV_D    = 32'b0001101??????????????????1010011;
    localparam [31:0] FSQRT_D   = 32'b010110100000?????????????1010011;
    localparam [31:0] FSGNJ_D   = 32'b0010001??????????000?????1010011;
    localparam [31:0] FSGNJN_D  = 32'b0010001??????????001?????1010011;
    localparam [31:0] FSGNJX_D  = 32'b0010001??????????010?????1010011;
    localparam [31:0] FMIN_D    = 32'b0010101??????????000?????1010011;
    localparam [31:0] FMAX_D    = 32'b0010101??????????001?????1010011;
    localparam [31:0] FCVT_W_D  = 32'b110000100000?????????????1010011;
    localparam [31:0] FCVT_WU_D = 32'b110000100001?????????????1010011;
    localparam [31:0] FCVT_D_W  = 32'b110100100000?????????????1010011;
    localparam [31:0] FCVT_D_WU = 32'b110100100001?????????????1010011;
    localparam [31:0] FEQ_D     = 32'b1010001??????????010?????1010011;
    localparam [31:0] FLT_D     = 32'b1010001??????????001?????1010011;
    localparam [31:0] FLE_D     = 32'b1010001??????????000?????1010011;
    localparam [31:0] FLASS_D   = 32'b111000100000?????001?????1010011;
    localparam [31:0] FCVT_S_D  = 32'b010000000001?????????????1010011;
    localparam [31:0] FCVT_D_S  = 32'b010000100000?????????????1010011;


    logic [6:0] opcode;
    logic [6:0] fn7;
    logic [4:0] opcode_trim;
    logic sp_legal;
    logic db_legal;
    //logic need_int_data;
    //logic write_int_data;
    //logic need_float_data;
    //logic write_float_data;
    logic instruction_is_float;
    ////////////////////////////////////////////////////
    //Implementation

    assign sp_legal = instruction inside {
        FLW, FSW, FMADD_S, FMSUB_S, FNMSUB_S, FNMADD_S, FADD_S, FSUB_S, FMUL_S,
        FDIV_S, FSQRT_S, FSGNJ_S, FSGNJN_S, FSGNJX_S, FMIN_S, FMAX_S, FCVT_W_S,
        FCVT_WU_S, FCVT_S_W, FCVT_S_WU, FMV_W_X, FMV_X_W, FEQ_S, FLT_S, FLE_S, FLASS_S
    };

    assign db_legal = instruction inside {
        FLD, FSD, FMADD_D, FMSUB_D, FNMSUB_D, FNMADD_D, FADD_D, FSUB_D, FMUL_D,
        FDIV_D, FSQRT_D, FSGNJ_D, FSGNJN_D, FSGNJX_D, FMIN_D, FMAX_D, FCVT_W_D,
        FCVT_WU_D, FCVT_D_W, FCVT_D_WU, FEQ_D, FLT_D, FLE_D, FLASS_D, FCVT_S_D, FCVT_D_S
    };

    //need to read from integer reg file
    assign need_int_data = instruction inside {
        FLW, FSW, FCVT_S_W, FCVT_S_WU, FMV_X_W,

        FLD, FSD, FCVT_D_W, FCVT_D_WU
    };

    assign need_float_data = instruction inside {
        FSW, FMADD_S, FMSUB_S, FNMSUB_S, FNMADD_S, FADD_S, FSUB_S, FMUL_S,
        FDIV_S, FSQRT_S, FSGNJ_S, FSGNJN_S, FSGNJX_S, FMIN_S, FMAX_S, FCVT_W_S,
        FCVT_WU_S, FMV_W_X, FEQ_S, FLT_S, FLE_S, FLASS_S,

        FSD, FMADD_D, FMSUB_D, FNMSUB_D, FNMADD_D, FADD_D, FSUB_D, FMUL_D,
        FDIV_D, FSQRT_D, FSGNJ_D, FSGNJN_D, FSGNJX_D, FMIN_D, FMAX_D, FCVT_W_D,
        FCVT_WU_D, FEQ_D, FLT_D, FLE_D, FLASS_D
    };

    //write back to integer reg file
    //assign write_int_data = instruction inside {
        //FCVT_W_S, FCVT_WU_S, FMV_X_W, FEQ_S, FLT_S, FLE_S, FLASS_S,

        //FCVT_W_D, FCVT_WU_D, FEQ_D, FLT_D, FLE_D, FLASS_D
    //};

    //assign write_float_data = instruction inside {
        //FLW, FMADD_S, FMSUB_S, FNMSUB_S, FNMADD_S, FADD_S, FSUB_S, FMUL_S,
        //FDIV_S, FSQRT_S, FSGNJ_S, FSGNJN_S, FSGNJX_S, FMIN_S, FMAX_S, FCVT_S_W, FCVT_S_WU, FMV_X_W,

        //FLD, FMADD_D, FMSUB_D, FNMSUB_D, FNMADD_D, FADD_D, FSUB_D, FMUL_D,
        //FDIV_D, FSQRT_D, FSGNJ_D, FSGNJN_D, FSGNJX_D, FMIN_D, FMAX_D, FCVT_D_W, FCVT_D_WU, FCVT_D_S, FCVT_S_D
    //};

    assign opcode = instruction[6:0];
    assign opcode_trim = opcode[6:2];
    assign fn7 = instruction[31:25];
    assign float_instruction = opcode_trim inside {FLD_T, FSD_T, FMADD_T, FMSUB_T, FNMSUB_T, FNMADD_T, FOP_T};//sp_legal | db_legal;
    assign write_int_data = (opcode_trim == FOP_T) & (fn7 inside {FCVT_WD, FCMP, FCLASS});
    assign write_float_data = float_instruction && !write_int_data && !(opcode_trim == FSD_T);

    assign accumulating_csrs = instruction inside {FMADD_D, FMSUB_D, FNMSUB_D, FNMADD_D,
        FMADD_D, FADD_D, FSUB_D, FMUL_D, FDIV_D, FSQRT_D, FMIN_D, FMAX_D, FCVT_S_D, FCVT_D_S,
        FEQ_D, FLT_D, FLE_D, FCVT_W_D, FCVT_WU_D
    };

endmodule
