/*
 * Copyright © 2017-2019 Eric Matthews,  Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Eric Matthews <ematthew@sfu.ca>
 */

module decode_and_issue

    import cva5_config::*;
    import riscv_types::*;
    import cva5_types::*;
    import csr_types::*;
    import opcodes::*;

    # (
        parameter cpu_config_t CONFIG = EXAMPLE_CONFIG
    )

    (
        input logic clk,
        input logic rst,

        //ID Management
        input logic pc_id_available,
        input decode_packet_t decode,
        output logic decode_advance,
        output exception_sources_t decode_exception_unit,

        //Renamer
        renamer_interface.decode renamer,

        input logic [MAX_NUM_UNITS-1:0] unit_needed,
        input logic [MAX_NUM_UNITS-1:0][REGFILE_READ_PORTS-1:0] unit_uses_rs,
        input logic [MAX_NUM_UNITS-1:0] unit_uses_rd,

        output logic decode_uses_rd,
        output rs_addr_t decode_rd_addr,
        output phys_addr_t decode_phys_rd_addr,
        output phys_addr_t decode_phys_rs_addr [REGFILE_READ_PORTS],
        output logic [$clog2(CONFIG.NUM_WB_GROUPS)-1:0] decode_rs_wb_group [REGFILE_READ_PORTS],

        output logic instruction_issued,
        output logic instruction_issued_with_rd,
        output issue_packet_t issue,
        output rs_addr_t issue_rs_addr [REGFILE_READ_PORTS],
        output phys_addr_t issue_phys_rs_addr [REGFILE_READ_PORTS],
        output logic [$clog2(CONFIG.NUM_WB_GROUPS)-1:0] issue_rd_wb_group,
        output logic issue_stage_ready,

        //Register File
        register_file_issue_interface.issue rf,

        output logic [31:0] constant_alu,

        unit_issue_interface.decode unit_issue [MAX_NUM_UNITS-1:0],

        input gc_outputs_t gc,
        input logic [1:0] current_privilege,

        exception_interface.unit exception
    );


    common_instruction_t decode_instruction;//rs1_addr, rs2_addr, fn3, fn7, rd_addr, upper/lower opcode

    logic decode_uses_rs [REGFILE_READ_PORTS];

    rs_addr_t decode_rs_addr [REGFILE_READ_PORTS];
    logic [$clog2(CONFIG.NUM_WB_GROUPS)-1:0] decode_wb_group;

    logic issue_hold;
    logic [REGFILE_READ_PORTS-1:0] operand_ready;
    logic [MAX_NUM_UNITS-1:0] unit_needed_issue_stage;
    logic [MAX_NUM_UNITS-1:0] issue_to;

    logic [$clog2(CONFIG.NUM_WB_GROUPS)-1:0] issue_rs_wb_group [REGFILE_READ_PORTS];
    logic issue_uses_rs [REGFILE_READ_PORTS];

    logic pre_issue_exception_pending;
    logic illegal_instruction_pattern;

    genvar i;
    ////////////////////////////////////////////////////
    //Implementation

    //Can move data into issue stage if:
    // there is no instruction currently in the issue stage, or
    // an instruction could issue (ignoring gc.fetch_flush)
    assign issue_stage_ready = (~issue.stage_valid) | (|issue_to);
    assign decode_advance = decode.valid & issue_stage_ready;

    //Instruction aliases
    assign decode_instruction = decode.instruction;
    always_comb begin
        decode_rs_addr = '{default: '0};
        decode_rs_addr[RS1] = decode_instruction.rs1_addr;
        decode_rs_addr[RS2] = decode_instruction.rs2_addr;
    end
    ////////////////////////////////////////////////////
    //Register File Support
    always_comb begin
        decode_uses_rd = |unit_uses_rd;
        decode_uses_rs = '{default: 0};
        for (int i = 0; i < MAX_NUM_UNITS; i++)
            for (int j = 0; j < REGFILE_READ_PORTS; j++)
                decode_uses_rs[j] |= unit_uses_rs[i][j];
    end

    ////////////////////////////////////////////////////
    //WB Group Determination
    localparam units_t [MAX_NUM_UNITS-1:0] WB_UNITS_TYPE_REP  = get_wb_units_type_representation(CONFIG.WB_GROUP);
    logic [CONFIG.NUM_WB_GROUPS-1:0] uses_wb_group;
    
    always_comb begin
        for (int i = 0; i < CONFIG.NUM_WB_GROUPS; i++)
            uses_wb_group[i] = |(unit_needed & WB_UNITS_TYPE_REP[i]);
    end

    one_hot_to_integer #(.C_WIDTH(CONFIG.NUM_WB_GROUPS))
    wb_group_one_hot_block (
        .one_hot (uses_wb_group),
        .int_out (decode_wb_group)
    );

    ////////////////////////////////////////////////////
    //Renamer Support
    assign renamer.rd_addr = decode_instruction.rd_addr;
    assign renamer.rs_addr = decode_rs_addr;
    assign renamer.uses_rd = decode_uses_rd;
    assign renamer.rd_wb_group = decode_wb_group;
    assign renamer.id = decode.id;

    ////////////////////////////////////////////////////
    //Decode ID Support
    assign decode_rd_addr = decode_instruction.rd_addr;
    assign decode_phys_rd_addr = renamer.phys_rd_addr;
    assign decode_phys_rs_addr = renamer.phys_rs_addr;
    assign decode_rs_wb_group = renamer.rs_wb_group;

    ////////////////////////////////////////////////////
    //Issue
    always_ff @(posedge clk) begin
        if (issue_stage_ready) begin
            issue.pc <= decode.pc;
            issue.instruction <= decode.instruction;
            issue.fetch_metadata <= decode.fetch_metadata;
            issue.fn3 <= decode_instruction.fn3;
            issue.opcode <= decode.instruction[6:0];
            issue_rs_addr <= decode_rs_addr;
            issue_phys_rs_addr <= renamer.phys_rs_addr;
            issue_rs_wb_group <= renamer.rs_wb_group;
            issue.rd_addr <= decode_instruction.rd_addr;
            issue.phys_rd_addr <= renamer.phys_rd_addr;
            issue_rd_wb_group <= decode_wb_group;
            issue.is_multicycle <= ~unit_needed[ALU_ID];
            issue.id <= decode.id;
            issue.exception_unit <= decode_exception_unit;
            issue_uses_rs <= decode_uses_rs;
            issue.uses_rd <= decode_uses_rd;
        end
    end

    always_ff @(posedge clk) begin
        if (issue_stage_ready)
            unit_needed_issue_stage <= unit_needed;
    end

    always_ff @(posedge clk) begin
        if (rst | gc.fetch_flush)
            issue.stage_valid <= 0;
        else if (issue_stage_ready)
            issue.stage_valid <= decode.valid;
    end

    ////////////////////////////////////////////////////
    //Issue Determination
    assign issue_hold = gc.issue_hold | pre_issue_exception_pending;

    generate for (i=0; i<REGFILE_READ_PORTS; i++)
        assign operand_ready[i] = ~rf.inuse[i] | (rf.inuse[i] & ~issue_uses_rs[i]);
    endgenerate

    ////////////////////////////////////////////////////
    //Unit EX signals
    generate for (i = 0; i < MAX_NUM_UNITS; i++) begin : gen_unit_issue_signals
        assign unit_issue[i].possible_issue = issue.stage_valid & unit_needed_issue_stage[i] & unit_issue[i].ready;
        assign issue_to[i] = unit_issue[i].possible_issue & (&operand_ready) & ~issue_hold;
        assign unit_issue[i].new_request = issue_to[i] & ~gc.fetch_flush;
        assign unit_issue[i].id = issue.id;
    end endgenerate

    assign instruction_issued = |issue_to & ~gc.fetch_flush;
    assign instruction_issued_with_rd = instruction_issued & issue.uses_rd;

    ////////////////////////////////////////////////////
    //Register File Issue Interface
    assign rf.phys_rs_addr = issue_phys_rs_addr;
    assign rf.phys_rd_addr = issue.phys_rd_addr;
    assign rf.rs_wb_group = issue_rs_wb_group;
    
    assign rf.single_cycle_or_flush = (instruction_issued_with_rd & |issue.rd_addr & ~issue.is_multicycle) | (issue.stage_valid & issue.uses_rd & |issue.rd_addr & gc.fetch_flush);
    
    ////////////////////////////////////////////////////
    //Constant ALU:
    //  provides LUI, AUIPC, JAL, JALR results for ALU
    //  provides PC+4 for BRANCH unit and ifence in GC unit
    always_ff @(posedge clk) begin
        if (issue_stage_ready)
            constant_alu <= ((decode_instruction.upper_opcode inside {LUI_T}) ? '0 : decode.pc) + ((decode_instruction.upper_opcode inside {LUI_T, AUIPC_T}) ? {decode.instruction[31:12], 12'b0} : 4); 
    end

    ////////////////////////////////////////////////////
    //Illegal Instruction check
    generate if (CONFIG.INCLUDE_M_MODE) begin : gen_decode_exceptions
    logic new_exception;
    exception_code_t ecode;
    exception_code_t ecall_code;

    //ECALL and EBREAK captured here, but seperated out when ecode is set
    assign illegal_instruction_pattern = ~|unit_needed;

    //TODO: Consider ways of parameterizing so that any exception generating unit
    //can be automatically added to this expression
    always_comb begin
        unique case (1'b1)
            unit_needed[LS_ID] : decode_exception_unit = LS_EXCEPTION;
            unit_needed[BR_ID] : decode_exception_unit = BR_EXCEPTION;
            default : decode_exception_unit = PRE_ISSUE_EXCEPTION;
        endcase
        if (~decode.fetch_metadata.ok)
            decode_exception_unit = PRE_ISSUE_EXCEPTION;
    end

    ////////////////////////////////////////////////////
    //ECALL/EBREAK
    //The type of call instruction is depedent on the current privilege level
    always_comb begin
        case (current_privilege)
            USER_PRIVILEGE : ecall_code = ECALL_U;
            SUPERVISOR_PRIVILEGE : ecall_code = ECALL_S;
            MACHINE_PRIVILEGE : ecall_code = ECALL_M;
            default : ecall_code = ECALL_U;
        endcase
    end

    always_ff @(posedge clk) begin
        if (issue_stage_ready) begin
            ecode <=
                    decode.instruction inside {ECALL} ? ecall_code :
                    decode.instruction inside {EBREAK} ? BREAK :
                    illegal_instruction_pattern ? ILLEGAL_INST :
                    decode.fetch_metadata.error_code; //(~decode.fetch_metadata.ok)
        end
    end

    ////////////////////////////////////////////////////
    //Exception generation (ecall/ebreak/illegal instruction/propagated fetch error)
    always_ff @(posedge clk) begin
        if (rst)
            pre_issue_exception_pending <= 0;
        else if (issue_stage_ready)
            pre_issue_exception_pending <= illegal_instruction_pattern | (~decode.fetch_metadata.ok);
    end

    assign new_exception = issue.stage_valid & pre_issue_exception_pending & ~(gc.issue_hold | gc.fetch_flush | exception.valid);

    always_ff @(posedge clk) begin
        if (rst)
            exception.valid <= 0;
        else
            exception.valid <= (exception.valid | new_exception) & ~exception.ack;
    end

    always_ff @(posedge clk) begin
        if (new_exception) begin
            exception.code <= ecode;
            exception.tval <= issue.instruction;
            exception.id <= issue.id;
        end
    end

    end endgenerate
    ////////////////////////////////////////////////////
    //End of Implementation
    ////////////////////////////////////////////////////

    ////////////////////////////////////////////////////
    //Assertions

endmodule
