/*
 * Copyright © 2023 Chris Keilbart, Lesley Shannon
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * Initial code developed under the supervision of Dr. Lesley Shannon,
 * Reconfigurable Computing Lab, Simon Fraser University.
 *
 * Author(s):
 *             Chris Keilbart <ckeilbar@sfu.ca>
 */

module q_lookup
    import fpu_types::*;

(
    input logic[2:0] d,
    input logic[6:0] ws,
    input logic[6:0] wc,
    output q_t q,
    output logic not_in_table //Only used for assertion
);

    logic[6:0] combined;
    assign combined = ws + wc;

    always_comb begin
        not_in_table = 0;
        //Table contents generated by genRadix4LUT.c
        unique case ({d, combined})
            10'b0001010100: q = NEG_TWO;
            10'b0001010101: q = NEG_TWO;
            10'b0001010110: q = NEG_TWO;
            10'b0001010111: q = NEG_TWO;
            10'b0001011000: q = NEG_TWO;
            10'b0001011001: q = NEG_TWO;
            10'b0001011010: q = NEG_TWO;
            10'b0001011011: q = NEG_TWO;
            10'b0001011100: q = NEG_TWO;
            10'b0001011101: q = NEG_TWO;
            10'b0001011110: q = NEG_TWO;
            10'b0001011111: q = NEG_TWO;
            10'b0001100000: q = NEG_TWO;
            10'b0001100001: q = NEG_TWO;
            10'b0001100010: q = NEG_TWO;
            10'b0001100011: q = NEG_TWO;
            10'b0001100100: q = NEG_TWO;
            10'b0001100101: q = NEG_TWO;
            10'b0001100110: q = NEG_TWO;
            10'b0001100111: q = NEG_TWO;
            10'b0001101000: q = NEG_TWO;
            10'b0001101001: q = NEG_TWO;
            10'b0001101010: q = NEG_TWO;
            10'b0001101011: q = NEG_TWO;
            10'b0001101100: q = NEG_TWO;
            10'b0001101101: q = NEG_TWO;
            10'b0001101110: q = NEG_TWO;
            10'b0001101111: q = NEG_TWO;
            10'b0001110000: q = NEG_TWO;
            10'b0001110001: q = NEG_TWO;
            10'b0001110010: q = NEG_TWO;
            10'b0001110011: q = NEG_ONE;
            10'b0001110100: q = NEG_ONE;
            10'b0001110101: q = NEG_ONE;
            10'b0001110110: q = NEG_ONE;
            10'b0001110111: q = NEG_ONE;
            10'b0001111000: q = NEG_ONE;
            10'b0001111001: q = NEG_ONE;
            10'b0001111010: q = NEG_ONE;
            10'b0001111011: q = NEG_ONE;
            10'b0001111100: q = ZERO;
            10'b0001111101: q = ZERO;
            10'b0001111110: q = ZERO;
            10'b0001111111: q = ZERO;
            10'b0000000000: q = ZERO;
            10'b0000000001: q = ZERO;
            10'b0000000010: q = ZERO;
            10'b0000000011: q = ZERO;
            10'b0000000100: q = POS_ONE;
            10'b0000000101: q = POS_ONE;
            10'b0000000110: q = POS_ONE;
            10'b0000000111: q = POS_ONE;
            10'b0000001000: q = POS_ONE;
            10'b0000001001: q = POS_ONE;
            10'b0000001010: q = POS_ONE;
            10'b0000001011: q = POS_ONE;
            10'b0000001100: q = POS_TWO;
            10'b0000001101: q = POS_TWO;
            10'b0000001110: q = POS_TWO;
            10'b0000001111: q = POS_TWO;
            10'b0000010000: q = POS_TWO;
            10'b0000010001: q = POS_TWO;
            10'b0000010010: q = POS_TWO;
            10'b0000010011: q = POS_TWO;
            10'b0000010100: q = POS_TWO;
            10'b0000010101: q = POS_TWO;
            10'b0000010110: q = POS_TWO;
            10'b0000010111: q = POS_TWO;
            10'b0000011000: q = POS_TWO;
            10'b0000011001: q = POS_TWO;
            10'b0000011010: q = POS_TWO;
            10'b0000011011: q = POS_TWO;
            10'b0000011100: q = POS_TWO;
            10'b0000011101: q = POS_TWO;
            10'b0000011110: q = POS_TWO;
            10'b0000011111: q = POS_TWO;
            10'b0000100000: q = POS_TWO;
            10'b0000100001: q = POS_TWO;
            10'b0000100010: q = POS_TWO;
            10'b0000100011: q = POS_TWO;
            10'b0000100100: q = POS_TWO;
            10'b0000100101: q = POS_TWO;
            10'b0000100110: q = POS_TWO;
            10'b0000100111: q = POS_TWO;
            10'b0000101000: q = POS_TWO;
            10'b0000101001: q = POS_TWO;
            10'b0000101010: q = POS_TWO;
            10'b0011010100: q = NEG_TWO;
            10'b0011010101: q = NEG_TWO;
            10'b0011010110: q = NEG_TWO;
            10'b0011010111: q = NEG_TWO;
            10'b0011011000: q = NEG_TWO;
            10'b0011011001: q = NEG_TWO;
            10'b0011011010: q = NEG_TWO;
            10'b0011011011: q = NEG_TWO;
            10'b0011011100: q = NEG_TWO;
            10'b0011011101: q = NEG_TWO;
            10'b0011011110: q = NEG_TWO;
            10'b0011011111: q = NEG_TWO;
            10'b0011100000: q = NEG_TWO;
            10'b0011100001: q = NEG_TWO;
            10'b0011100010: q = NEG_TWO;
            10'b0011100011: q = NEG_TWO;
            10'b0011100100: q = NEG_TWO;
            10'b0011100101: q = NEG_TWO;
            10'b0011100110: q = NEG_TWO;
            10'b0011100111: q = NEG_TWO;
            10'b0011101000: q = NEG_TWO;
            10'b0011101001: q = NEG_TWO;
            10'b0011101010: q = NEG_TWO;
            10'b0011101011: q = NEG_TWO;
            10'b0011101100: q = NEG_TWO;
            10'b0011101101: q = NEG_TWO;
            10'b0011101110: q = NEG_TWO;
            10'b0011101111: q = NEG_TWO;
            10'b0011110000: q = NEG_TWO;
            10'b0011110001: q = NEG_ONE;
            10'b0011110010: q = NEG_ONE;
            10'b0011110011: q = NEG_ONE;
            10'b0011110100: q = NEG_ONE;
            10'b0011110101: q = NEG_ONE;
            10'b0011110110: q = NEG_ONE;
            10'b0011110111: q = NEG_ONE;
            10'b0011111000: q = NEG_ONE;
            10'b0011111001: q = NEG_ONE;
            10'b0011111010: q = ZERO;
            10'b0011111011: q = ZERO;
            10'b0011111100: q = ZERO;
            10'b0011111101: q = ZERO;
            10'b0011111110: q = ZERO;
            10'b0011111111: q = ZERO;
            10'b0010000000: q = ZERO;
            10'b0010000001: q = ZERO;
            10'b0010000010: q = ZERO;
            10'b0010000011: q = ZERO;
            10'b0010000100: q = POS_ONE;
            10'b0010000101: q = POS_ONE;
            10'b0010000110: q = POS_ONE;
            10'b0010000111: q = POS_ONE;
            10'b0010001000: q = POS_ONE;
            10'b0010001001: q = POS_ONE;
            10'b0010001010: q = POS_ONE;
            10'b0010001011: q = POS_ONE;
            10'b0010001100: q = POS_ONE;
            10'b0010001101: q = POS_ONE;
            10'b0010001110: q = POS_TWO;
            10'b0010001111: q = POS_TWO;
            10'b0010010000: q = POS_TWO;
            10'b0010010001: q = POS_TWO;
            10'b0010010010: q = POS_TWO;
            10'b0010010011: q = POS_TWO;
            10'b0010010100: q = POS_TWO;
            10'b0010010101: q = POS_TWO;
            10'b0010010110: q = POS_TWO;
            10'b0010010111: q = POS_TWO;
            10'b0010011000: q = POS_TWO;
            10'b0010011001: q = POS_TWO;
            10'b0010011010: q = POS_TWO;
            10'b0010011011: q = POS_TWO;
            10'b0010011100: q = POS_TWO;
            10'b0010011101: q = POS_TWO;
            10'b0010011110: q = POS_TWO;
            10'b0010011111: q = POS_TWO;
            10'b0010100000: q = POS_TWO;
            10'b0010100001: q = POS_TWO;
            10'b0010100010: q = POS_TWO;
            10'b0010100011: q = POS_TWO;
            10'b0010100100: q = POS_TWO;
            10'b0010100101: q = POS_TWO;
            10'b0010100110: q = POS_TWO;
            10'b0010100111: q = POS_TWO;
            10'b0010101000: q = POS_TWO;
            10'b0010101001: q = POS_TWO;
            10'b0010101010: q = POS_TWO;
            10'b0101010100: q = NEG_TWO;
            10'b0101010101: q = NEG_TWO;
            10'b0101010110: q = NEG_TWO;
            10'b0101010111: q = NEG_TWO;
            10'b0101011000: q = NEG_TWO;
            10'b0101011001: q = NEG_TWO;
            10'b0101011010: q = NEG_TWO;
            10'b0101011011: q = NEG_TWO;
            10'b0101011100: q = NEG_TWO;
            10'b0101011101: q = NEG_TWO;
            10'b0101011110: q = NEG_TWO;
            10'b0101011111: q = NEG_TWO;
            10'b0101100000: q = NEG_TWO;
            10'b0101100001: q = NEG_TWO;
            10'b0101100010: q = NEG_TWO;
            10'b0101100011: q = NEG_TWO;
            10'b0101100100: q = NEG_TWO;
            10'b0101100101: q = NEG_TWO;
            10'b0101100110: q = NEG_TWO;
            10'b0101100111: q = NEG_TWO;
            10'b0101101000: q = NEG_TWO;
            10'b0101101001: q = NEG_TWO;
            10'b0101101010: q = NEG_TWO;
            10'b0101101011: q = NEG_TWO;
            10'b0101101100: q = NEG_TWO;
            10'b0101101101: q = NEG_TWO;
            10'b0101101110: q = NEG_TWO;
            10'b0101101111: q = NEG_TWO;
            10'b0101110000: q = NEG_ONE;
            10'b0101110001: q = NEG_ONE;
            10'b0101110010: q = NEG_ONE;
            10'b0101110011: q = NEG_ONE;
            10'b0101110100: q = NEG_ONE;
            10'b0101110101: q = NEG_ONE;
            10'b0101110110: q = NEG_ONE;
            10'b0101110111: q = NEG_ONE;
            10'b0101111000: q = NEG_ONE;
            10'b0101111001: q = NEG_ONE;
            10'b0101111010: q = ZERO;
            10'b0101111011: q = ZERO;
            10'b0101111100: q = ZERO;
            10'b0101111101: q = ZERO;
            10'b0101111110: q = ZERO;
            10'b0101111111: q = ZERO;
            10'b0100000000: q = ZERO;
            10'b0100000001: q = ZERO;
            10'b0100000010: q = ZERO;
            10'b0100000011: q = ZERO;
            10'b0100000100: q = POS_ONE;
            10'b0100000101: q = POS_ONE;
            10'b0100000110: q = POS_ONE;
            10'b0100000111: q = POS_ONE;
            10'b0100001000: q = POS_ONE;
            10'b0100001001: q = POS_ONE;
            10'b0100001010: q = POS_ONE;
            10'b0100001011: q = POS_ONE;
            10'b0100001100: q = POS_ONE;
            10'b0100001101: q = POS_ONE;
            10'b0100001110: q = POS_ONE;
            10'b0100001111: q = POS_TWO;
            10'b0100010000: q = POS_TWO;
            10'b0100010001: q = POS_TWO;
            10'b0100010010: q = POS_TWO;
            10'b0100010011: q = POS_TWO;
            10'b0100010100: q = POS_TWO;
            10'b0100010101: q = POS_TWO;
            10'b0100010110: q = POS_TWO;
            10'b0100010111: q = POS_TWO;
            10'b0100011000: q = POS_TWO;
            10'b0100011001: q = POS_TWO;
            10'b0100011010: q = POS_TWO;
            10'b0100011011: q = POS_TWO;
            10'b0100011100: q = POS_TWO;
            10'b0100011101: q = POS_TWO;
            10'b0100011110: q = POS_TWO;
            10'b0100011111: q = POS_TWO;
            10'b0100100000: q = POS_TWO;
            10'b0100100001: q = POS_TWO;
            10'b0100100010: q = POS_TWO;
            10'b0100100011: q = POS_TWO;
            10'b0100100100: q = POS_TWO;
            10'b0100100101: q = POS_TWO;
            10'b0100100110: q = POS_TWO;
            10'b0100100111: q = POS_TWO;
            10'b0100101000: q = POS_TWO;
            10'b0100101001: q = POS_TWO;
            10'b0100101010: q = POS_TWO;
            10'b0111010100: q = NEG_TWO;
            10'b0111010101: q = NEG_TWO;
            10'b0111010110: q = NEG_TWO;
            10'b0111010111: q = NEG_TWO;
            10'b0111011000: q = NEG_TWO;
            10'b0111011001: q = NEG_TWO;
            10'b0111011010: q = NEG_TWO;
            10'b0111011011: q = NEG_TWO;
            10'b0111011100: q = NEG_TWO;
            10'b0111011101: q = NEG_TWO;
            10'b0111011110: q = NEG_TWO;
            10'b0111011111: q = NEG_TWO;
            10'b0111100000: q = NEG_TWO;
            10'b0111100001: q = NEG_TWO;
            10'b0111100010: q = NEG_TWO;
            10'b0111100011: q = NEG_TWO;
            10'b0111100100: q = NEG_TWO;
            10'b0111100101: q = NEG_TWO;
            10'b0111100110: q = NEG_TWO;
            10'b0111100111: q = NEG_TWO;
            10'b0111101000: q = NEG_TWO;
            10'b0111101001: q = NEG_TWO;
            10'b0111101010: q = NEG_TWO;
            10'b0111101011: q = NEG_TWO;
            10'b0111101100: q = NEG_TWO;
            10'b0111101101: q = NEG_TWO;
            10'b0111101110: q = NEG_ONE;
            10'b0111101111: q = NEG_ONE;
            10'b0111110000: q = NEG_ONE;
            10'b0111110001: q = NEG_ONE;
            10'b0111110010: q = NEG_ONE;
            10'b0111110011: q = NEG_ONE;
            10'b0111110100: q = NEG_ONE;
            10'b0111110101: q = NEG_ONE;
            10'b0111110110: q = NEG_ONE;
            10'b0111110111: q = NEG_ONE;
            10'b0111111000: q = NEG_ONE;
            10'b0111111001: q = NEG_ONE;
            10'b0111111010: q = ZERO;
            10'b0111111011: q = ZERO;
            10'b0111111100: q = ZERO;
            10'b0111111101: q = ZERO;
            10'b0111111110: q = ZERO;
            10'b0111111111: q = ZERO;
            10'b0110000000: q = ZERO;
            10'b0110000001: q = ZERO;
            10'b0110000010: q = ZERO;
            10'b0110000011: q = ZERO;
            10'b0110000100: q = POS_ONE;
            10'b0110000101: q = POS_ONE;
            10'b0110000110: q = POS_ONE;
            10'b0110000111: q = POS_ONE;
            10'b0110001000: q = POS_ONE;
            10'b0110001001: q = POS_ONE;
            10'b0110001010: q = POS_ONE;
            10'b0110001011: q = POS_ONE;
            10'b0110001100: q = POS_ONE;
            10'b0110001101: q = POS_ONE;
            10'b0110001110: q = POS_ONE;
            10'b0110001111: q = POS_ONE;
            10'b0110010000: q = POS_TWO;
            10'b0110010001: q = POS_TWO;
            10'b0110010010: q = POS_TWO;
            10'b0110010011: q = POS_TWO;
            10'b0110010100: q = POS_TWO;
            10'b0110010101: q = POS_TWO;
            10'b0110010110: q = POS_TWO;
            10'b0110010111: q = POS_TWO;
            10'b0110011000: q = POS_TWO;
            10'b0110011001: q = POS_TWO;
            10'b0110011010: q = POS_TWO;
            10'b0110011011: q = POS_TWO;
            10'b0110011100: q = POS_TWO;
            10'b0110011101: q = POS_TWO;
            10'b0110011110: q = POS_TWO;
            10'b0110011111: q = POS_TWO;
            10'b0110100000: q = POS_TWO;
            10'b0110100001: q = POS_TWO;
            10'b0110100010: q = POS_TWO;
            10'b0110100011: q = POS_TWO;
            10'b0110100100: q = POS_TWO;
            10'b0110100101: q = POS_TWO;
            10'b0110100110: q = POS_TWO;
            10'b0110100111: q = POS_TWO;
            10'b0110101000: q = POS_TWO;
            10'b0110101001: q = POS_TWO;
            10'b0110101010: q = POS_TWO;
            10'b1001010100: q = NEG_TWO;
            10'b1001010101: q = NEG_TWO;
            10'b1001010110: q = NEG_TWO;
            10'b1001010111: q = NEG_TWO;
            10'b1001011000: q = NEG_TWO;
            10'b1001011001: q = NEG_TWO;
            10'b1001011010: q = NEG_TWO;
            10'b1001011011: q = NEG_TWO;
            10'b1001011100: q = NEG_TWO;
            10'b1001011101: q = NEG_TWO;
            10'b1001011110: q = NEG_TWO;
            10'b1001011111: q = NEG_TWO;
            10'b1001100000: q = NEG_TWO;
            10'b1001100001: q = NEG_TWO;
            10'b1001100010: q = NEG_TWO;
            10'b1001100011: q = NEG_TWO;
            10'b1001100100: q = NEG_TWO;
            10'b1001100101: q = NEG_TWO;
            10'b1001100110: q = NEG_TWO;
            10'b1001100111: q = NEG_TWO;
            10'b1001101000: q = NEG_TWO;
            10'b1001101001: q = NEG_TWO;
            10'b1001101010: q = NEG_TWO;
            10'b1001101011: q = NEG_TWO;
            10'b1001101100: q = NEG_ONE;
            10'b1001101101: q = NEG_ONE;
            10'b1001101110: q = NEG_ONE;
            10'b1001101111: q = NEG_ONE;
            10'b1001110000: q = NEG_ONE;
            10'b1001110001: q = NEG_ONE;
            10'b1001110010: q = NEG_ONE;
            10'b1001110011: q = NEG_ONE;
            10'b1001110100: q = NEG_ONE;
            10'b1001110101: q = NEG_ONE;
            10'b1001110110: q = NEG_ONE;
            10'b1001110111: q = NEG_ONE;
            10'b1001111000: q = ZERO;
            10'b1001111001: q = ZERO;
            10'b1001111010: q = ZERO;
            10'b1001111011: q = ZERO;
            10'b1001111100: q = ZERO;
            10'b1001111101: q = ZERO;
            10'b1001111110: q = ZERO;
            10'b1001111111: q = ZERO;
            10'b1000000000: q = ZERO;
            10'b1000000001: q = ZERO;
            10'b1000000010: q = ZERO;
            10'b1000000011: q = ZERO;
            10'b1000000100: q = ZERO;
            10'b1000000101: q = ZERO;
            10'b1000000110: q = POS_ONE;
            10'b1000000111: q = POS_ONE;
            10'b1000001000: q = POS_ONE;
            10'b1000001001: q = POS_ONE;
            10'b1000001010: q = POS_ONE;
            10'b1000001011: q = POS_ONE;
            10'b1000001100: q = POS_ONE;
            10'b1000001101: q = POS_ONE;
            10'b1000001110: q = POS_ONE;
            10'b1000001111: q = POS_ONE;
            10'b1000010000: q = POS_ONE;
            10'b1000010001: q = POS_ONE;
            10'b1000010010: q = POS_TWO;
            10'b1000010011: q = POS_TWO;
            10'b1000010100: q = POS_TWO;
            10'b1000010101: q = POS_TWO;
            10'b1000010110: q = POS_TWO;
            10'b1000010111: q = POS_TWO;
            10'b1000011000: q = POS_TWO;
            10'b1000011001: q = POS_TWO;
            10'b1000011010: q = POS_TWO;
            10'b1000011011: q = POS_TWO;
            10'b1000011100: q = POS_TWO;
            10'b1000011101: q = POS_TWO;
            10'b1000011110: q = POS_TWO;
            10'b1000011111: q = POS_TWO;
            10'b1000100000: q = POS_TWO;
            10'b1000100001: q = POS_TWO;
            10'b1000100010: q = POS_TWO;
            10'b1000100011: q = POS_TWO;
            10'b1000100100: q = POS_TWO;
            10'b1000100101: q = POS_TWO;
            10'b1000100110: q = POS_TWO;
            10'b1000100111: q = POS_TWO;
            10'b1000101000: q = POS_TWO;
            10'b1000101001: q = POS_TWO;
            10'b1000101010: q = POS_TWO;
            10'b1011010100: q = NEG_TWO;
            10'b1011010101: q = NEG_TWO;
            10'b1011010110: q = NEG_TWO;
            10'b1011010111: q = NEG_TWO;
            10'b1011011000: q = NEG_TWO;
            10'b1011011001: q = NEG_TWO;
            10'b1011011010: q = NEG_TWO;
            10'b1011011011: q = NEG_TWO;
            10'b1011011100: q = NEG_TWO;
            10'b1011011101: q = NEG_TWO;
            10'b1011011110: q = NEG_TWO;
            10'b1011011111: q = NEG_TWO;
            10'b1011100000: q = NEG_TWO;
            10'b1011100001: q = NEG_TWO;
            10'b1011100010: q = NEG_TWO;
            10'b1011100011: q = NEG_TWO;
            10'b1011100100: q = NEG_TWO;
            10'b1011100101: q = NEG_TWO;
            10'b1011100110: q = NEG_TWO;
            10'b1011100111: q = NEG_TWO;
            10'b1011101000: q = NEG_TWO;
            10'b1011101001: q = NEG_TWO;
            10'b1011101010: q = NEG_TWO;
            10'b1011101011: q = NEG_TWO;
            10'b1011101100: q = NEG_ONE;
            10'b1011101101: q = NEG_ONE;
            10'b1011101110: q = NEG_ONE;
            10'b1011101111: q = NEG_ONE;
            10'b1011110000: q = NEG_ONE;
            10'b1011110001: q = NEG_ONE;
            10'b1011110010: q = NEG_ONE;
            10'b1011110011: q = NEG_ONE;
            10'b1011110100: q = NEG_ONE;
            10'b1011110101: q = NEG_ONE;
            10'b1011110110: q = NEG_ONE;
            10'b1011110111: q = NEG_ONE;
            10'b1011111000: q = ZERO;
            10'b1011111001: q = ZERO;
            10'b1011111010: q = ZERO;
            10'b1011111011: q = ZERO;
            10'b1011111100: q = ZERO;
            10'b1011111101: q = ZERO;
            10'b1011111110: q = ZERO;
            10'b1011111111: q = ZERO;
            10'b1010000000: q = ZERO;
            10'b1010000001: q = ZERO;
            10'b1010000010: q = ZERO;
            10'b1010000011: q = ZERO;
            10'b1010000100: q = ZERO;
            10'b1010000101: q = ZERO;
            10'b1010000110: q = POS_ONE;
            10'b1010000111: q = POS_ONE;
            10'b1010001000: q = POS_ONE;
            10'b1010001001: q = POS_ONE;
            10'b1010001010: q = POS_ONE;
            10'b1010001011: q = POS_ONE;
            10'b1010001100: q = POS_ONE;
            10'b1010001101: q = POS_ONE;
            10'b1010001110: q = POS_ONE;
            10'b1010001111: q = POS_ONE;
            10'b1010010000: q = POS_ONE;
            10'b1010010001: q = POS_ONE;
            10'b1010010010: q = POS_ONE;
            10'b1010010011: q = POS_ONE;
            10'b1010010100: q = POS_TWO;
            10'b1010010101: q = POS_TWO;
            10'b1010010110: q = POS_TWO;
            10'b1010010111: q = POS_TWO;
            10'b1010011000: q = POS_TWO;
            10'b1010011001: q = POS_TWO;
            10'b1010011010: q = POS_TWO;
            10'b1010011011: q = POS_TWO;
            10'b1010011100: q = POS_TWO;
            10'b1010011101: q = POS_TWO;
            10'b1010011110: q = POS_TWO;
            10'b1010011111: q = POS_TWO;
            10'b1010100000: q = POS_TWO;
            10'b1010100001: q = POS_TWO;
            10'b1010100010: q = POS_TWO;
            10'b1010100011: q = POS_TWO;
            10'b1010100100: q = POS_TWO;
            10'b1010100101: q = POS_TWO;
            10'b1010100110: q = POS_TWO;
            10'b1010100111: q = POS_TWO;
            10'b1010101000: q = POS_TWO;
            10'b1010101001: q = POS_TWO;
            10'b1010101010: q = POS_TWO;
            10'b1101010100: q = NEG_TWO;
            10'b1101010101: q = NEG_TWO;
            10'b1101010110: q = NEG_TWO;
            10'b1101010111: q = NEG_TWO;
            10'b1101011000: q = NEG_TWO;
            10'b1101011001: q = NEG_TWO;
            10'b1101011010: q = NEG_TWO;
            10'b1101011011: q = NEG_TWO;
            10'b1101011100: q = NEG_TWO;
            10'b1101011101: q = NEG_TWO;
            10'b1101011110: q = NEG_TWO;
            10'b1101011111: q = NEG_TWO;
            10'b1101100000: q = NEG_TWO;
            10'b1101100001: q = NEG_TWO;
            10'b1101100010: q = NEG_TWO;
            10'b1101100011: q = NEG_TWO;
            10'b1101100100: q = NEG_TWO;
            10'b1101100101: q = NEG_TWO;
            10'b1101100110: q = NEG_TWO;
            10'b1101100111: q = NEG_TWO;
            10'b1101101000: q = NEG_TWO;
            10'b1101101001: q = NEG_TWO;
            10'b1101101010: q = NEG_ONE;
            10'b1101101011: q = NEG_ONE;
            10'b1101101100: q = NEG_ONE;
            10'b1101101101: q = NEG_ONE;
            10'b1101101110: q = NEG_ONE;
            10'b1101101111: q = NEG_ONE;
            10'b1101110000: q = NEG_ONE;
            10'b1101110001: q = NEG_ONE;
            10'b1101110010: q = NEG_ONE;
            10'b1101110011: q = NEG_ONE;
            10'b1101110100: q = NEG_ONE;
            10'b1101110101: q = NEG_ONE;
            10'b1101110110: q = NEG_ONE;
            10'b1101110111: q = NEG_ONE;
            10'b1101111000: q = ZERO;
            10'b1101111001: q = ZERO;
            10'b1101111010: q = ZERO;
            10'b1101111011: q = ZERO;
            10'b1101111100: q = ZERO;
            10'b1101111101: q = ZERO;
            10'b1101111110: q = ZERO;
            10'b1101111111: q = ZERO;
            10'b1100000000: q = ZERO;
            10'b1100000001: q = ZERO;
            10'b1100000010: q = ZERO;
            10'b1100000011: q = ZERO;
            10'b1100000100: q = ZERO;
            10'b1100000101: q = ZERO;
            10'b1100000110: q = ZERO;
            10'b1100000111: q = ZERO;
            10'b1100001000: q = POS_ONE;
            10'b1100001001: q = POS_ONE;
            10'b1100001010: q = POS_ONE;
            10'b1100001011: q = POS_ONE;
            10'b1100001100: q = POS_ONE;
            10'b1100001101: q = POS_ONE;
            10'b1100001110: q = POS_ONE;
            10'b1100001111: q = POS_ONE;
            10'b1100010000: q = POS_ONE;
            10'b1100010001: q = POS_ONE;
            10'b1100010010: q = POS_ONE;
            10'b1100010011: q = POS_ONE;
            10'b1100010100: q = POS_TWO;
            10'b1100010101: q = POS_TWO;
            10'b1100010110: q = POS_TWO;
            10'b1100010111: q = POS_TWO;
            10'b1100011000: q = POS_TWO;
            10'b1100011001: q = POS_TWO;
            10'b1100011010: q = POS_TWO;
            10'b1100011011: q = POS_TWO;
            10'b1100011100: q = POS_TWO;
            10'b1100011101: q = POS_TWO;
            10'b1100011110: q = POS_TWO;
            10'b1100011111: q = POS_TWO;
            10'b1100100000: q = POS_TWO;
            10'b1100100001: q = POS_TWO;
            10'b1100100010: q = POS_TWO;
            10'b1100100011: q = POS_TWO;
            10'b1100100100: q = POS_TWO;
            10'b1100100101: q = POS_TWO;
            10'b1100100110: q = POS_TWO;
            10'b1100100111: q = POS_TWO;
            10'b1100101000: q = POS_TWO;
            10'b1100101001: q = POS_TWO;
            10'b1100101010: q = POS_TWO;
            10'b1111010100: q = NEG_TWO;
            10'b1111010101: q = NEG_TWO;
            10'b1111010110: q = NEG_TWO;
            10'b1111010111: q = NEG_TWO;
            10'b1111011000: q = NEG_TWO;
            10'b1111011001: q = NEG_TWO;
            10'b1111011010: q = NEG_TWO;
            10'b1111011011: q = NEG_TWO;
            10'b1111011100: q = NEG_TWO;
            10'b1111011101: q = NEG_TWO;
            10'b1111011110: q = NEG_TWO;
            10'b1111011111: q = NEG_TWO;
            10'b1111100000: q = NEG_TWO;
            10'b1111100001: q = NEG_TWO;
            10'b1111100010: q = NEG_TWO;
            10'b1111100011: q = NEG_TWO;
            10'b1111100100: q = NEG_TWO;
            10'b1111100101: q = NEG_TWO;
            10'b1111100110: q = NEG_TWO;
            10'b1111100111: q = NEG_TWO;
            10'b1111101000: q = NEG_ONE;
            10'b1111101001: q = NEG_ONE;
            10'b1111101010: q = NEG_ONE;
            10'b1111101011: q = NEG_ONE;
            10'b1111101100: q = NEG_ONE;
            10'b1111101101: q = NEG_ONE;
            10'b1111101110: q = NEG_ONE;
            10'b1111101111: q = NEG_ONE;
            10'b1111110000: q = NEG_ONE;
            10'b1111110001: q = NEG_ONE;
            10'b1111110010: q = NEG_ONE;
            10'b1111110011: q = NEG_ONE;
            10'b1111110100: q = NEG_ONE;
            10'b1111110101: q = NEG_ONE;
            10'b1111110110: q = NEG_ONE;
            10'b1111110111: q = NEG_ONE;
            10'b1111111000: q = ZERO;
            10'b1111111001: q = ZERO;
            10'b1111111010: q = ZERO;
            10'b1111111011: q = ZERO;
            10'b1111111100: q = ZERO;
            10'b1111111101: q = ZERO;
            10'b1111111110: q = ZERO;
            10'b1111111111: q = ZERO;
            10'b1110000000: q = ZERO;
            10'b1110000001: q = ZERO;
            10'b1110000010: q = ZERO;
            10'b1110000011: q = ZERO;
            10'b1110000100: q = ZERO;
            10'b1110000101: q = ZERO;
            10'b1110000110: q = ZERO;
            10'b1110000111: q = ZERO;
            10'b1110001000: q = POS_ONE;
            10'b1110001001: q = POS_ONE;
            10'b1110001010: q = POS_ONE;
            10'b1110001011: q = POS_ONE;
            10'b1110001100: q = POS_ONE;
            10'b1110001101: q = POS_ONE;
            10'b1110001110: q = POS_ONE;
            10'b1110001111: q = POS_ONE;
            10'b1110010000: q = POS_ONE;
            10'b1110010001: q = POS_ONE;
            10'b1110010010: q = POS_ONE;
            10'b1110010011: q = POS_ONE;
            10'b1110010100: q = POS_ONE;
            10'b1110010101: q = POS_ONE;
            10'b1110010110: q = POS_ONE;
            10'b1110010111: q = POS_ONE;
            10'b1110011000: q = POS_TWO;
            10'b1110011001: q = POS_TWO;
            10'b1110011010: q = POS_TWO;
            10'b1110011011: q = POS_TWO;
            10'b1110011100: q = POS_TWO;
            10'b1110011101: q = POS_TWO;
            10'b1110011110: q = POS_TWO;
            10'b1110011111: q = POS_TWO;
            10'b1110100000: q = POS_TWO;
            10'b1110100001: q = POS_TWO;
            10'b1110100010: q = POS_TWO;
            10'b1110100011: q = POS_TWO;
            10'b1110100100: q = POS_TWO;
            10'b1110100101: q = POS_TWO;
            10'b1110100110: q = POS_TWO;
            10'b1110100111: q = POS_TWO;
            10'b1110101000: q = POS_TWO;
            10'b1110101001: q = POS_TWO;
            10'b1110101010: q = POS_TWO;
            default: begin //This should never be reached
                q = q_t'(3'bXXX); //This prevents the tool from creating potentially costly default behaviour
                not_in_table = 1;
            end
        endcase
    end

endmodule